* Qucs 2.0.0 /home/arficx/Desktop/circuits/LNA/qucs-sims/LNA-sim.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 2.0.0  /home/arficx/Desktop/circuits/LNA/qucs-sims/LNA-sim.sch

** sch_path: /home/arficx/Desktop/circuits/LNA/LNA-spice.sch
.subckt LNA-spice b g d s
XM1 d g s b sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends
.end

.LIB "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.PARAM vg = 900m

Xnfet_01v8_lvt 0 _net0 _net1 0 LNA-spice
EPr1 Pr1 0 _net0 0 1.0
RPr1Pr1 Pr1 0 1E8
RPr1_net0 _net0 0 1E8
Vid _net3 _net1 DC 0
V2 _net3 0 DC 1
vg _net0 0 DC {VG}
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz


save all

save @m.Xnfet_01v8_lvt.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.Xnfet_01v8_lvt.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]


dc vg -0.2 1.8 1m

let idn=@m.Xnfet_01v8_lvt.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
let gm=@m.Xnfet_01v8_lvt.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]

let gmoverid=gm/idn


write LNA-sim_custom.txt V(Pr1) Vid#branch idn gm gmoverid
destroy all
reset
exit
.endc
.END
