** sch_path: /home/engg/Desktop/IC Design/gmid_char/PMOS_Charac/pmos_gmid.sch
**.subckt pmos_gmid
XM1 net2 net1 GND GND sky130_fd_pr__pfet_01v8 L='length' W='width' nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 GND net1 0.9
V2 GND net2 0.9
**** begin user architecture code



.include init.txt
.include pmos_params.txt

.param length = 0.3
.param width = 1






**** end user architecture code
**.ends
.GLOBAL GND
.end
