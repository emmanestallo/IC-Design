** sch_path: /home/engg/Desktop/IC Design/test.sch
**.subckt test
V1 net1 GND 1
V2 net2 GND 1
XM1 net1 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1

.control
save all

save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]

dc v2 0 1 1m

let gm = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let id = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
let gds = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let cgg = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
let vdsat = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]

let gain = gm/gds
let ft = gm/(2*3.1415*cgg)
let gmoverid = gm/id

plot gain
plot ft
plot gmoverid
plot id
plot vdsat

wrdata gain.txt gain
wrdata ft.txt ft
wrdata gmoverid.txt gmoverid
wrdata id.txt id

.endc




**** end user architecture code
**.ends
.GLOBAL GND
.end
