* Qucs 2.0.0 /home/arficx/Desktop/circuits/LNA/s-param.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 2.0.0  /home/arficx/Desktop/circuits/LNA/s-param.sch
.LIB "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
