** sch_path: /home/engg/Desktop/IC Design/RF/RLC_Networks/parallel_rlc_tank.sch
**.subckt parallel_rlc_tank
L1 out GND 1n m=1
R1 out GND 1k m=1
C1 out GND 1p m=1
I0 out GND 10m AC 1
**** begin user architecture code



.control
save all
ac dec 10 1 100T
plot db(v(out))


.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
