** sch_path: /home/engg/Desktop/IC Design/gmid_char/test.sch
**.subckt test
V1 net1 GND 0.9
V2 net2 GND 0.9
XM1 net1 net2 GND GND sky130_fd_pr__nfet_01v8 L=length W=width nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1

.param length = 0.4
.param width = 1

.control
save all

save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8[id]
save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
save @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
save @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
save @m.xm1.msky130_fd_pr__nfet_01v8[vgs]

dc v2 0 1 1m

let gm = @m.xm1.msky130_fd_pr__nfet_01v8[gm]
let id = @m.xm1.msky130_fd_pr__nfet_01v8[id]
let gds = @m.xm1.msky130_fd_pr__nfet_01v8[gds]
let cgg = @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
let vdsat = @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
let vgs = @m.xm1.msky130_fd_pr__nfet_01v8[vgs]

let gmro = gm/gds
let ft = gm/(2*pi*cgg)
let gmoverid = gm/id

wrdata gmro.txt gmro
wrdata ft.txt ft
wrdata gmoverid.txt gmoverid
wrdata id.txt id
wrdata vdsat.txt vdsat
wrdata vgs.txt vgs

.endc




**** end user architecture code
**.ends
.GLOBAL GND
.end
