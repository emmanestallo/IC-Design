** sch_path: /home/emman/Desktop/IC-Design/BandgapReference/BGR_char.sch
**.subckt BGR_char
XM1 net1 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.6 W=11.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 net1 GND 0.9
**** begin user architecture code


.include init.txt

.control
save all

save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8[id]
save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
save @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
save @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
save @m.xm1.msky130_fd_pr__nfet_01v8[vgs]

dc v1 0 1 1m

let gm = @m.xm1.msky130_fd_pr__nfet_01v8[gm]
let id = @m.xm1.msky130_fd_pr__nfet_01v8[id]
let gds = @m.xm1.msky130_fd_pr__nfet_01v8[gds]
let cgg = @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
let vdsat = @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
let vgs = @m.xm1.msky130_fd_pr__nfet_01v8[vgs]

let gmro = gm/gds
let ft = gm/(2*pi*cgg)
let gmoverid = gm/id

.endc




**** end user architecture code
**.ends
.GLOBAL GND
.end
